/*
   Author: Ovidiu Plugariu
   Description: This is a test for the LZ77 sliding algorithm used in GZIP.  
*/
`include "gzip_pkg.sv"
import gzip_pkg::*;

module lz77_test();













endmodule
