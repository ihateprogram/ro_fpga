// This file has the 5 bit Huffman codes for Statis Distance Huffman Tree

`ifndef __huffman_dist_table__
`define __huffman_dist_table__

`define DIST_CODE0     5'd0   
`define DIST_CODE1     5'd1
`define DIST_CODE2     5'd2
`define DIST_CODE3     5'd3
`define DIST_CODE4     5'd4
`define DIST_CODE5     5'd5
`define DIST_CODE6     5'd6
`define DIST_CODE7     5'd7
`define DIST_CODE8     5'd8
`define DIST_CODE9     5'd9
`define DIST_CODE10    5'd10
`define DIST_CODE11    5'd11
`define DIST_CODE12    5'd12
`define DIST_CODE13    5'd13
`define DIST_CODE14    5'd14
`define DIST_CODE15    5'd15
`define DIST_CODE16    5'd16
`define DIST_CODE17    5'd17
`define DIST_CODE18    5'd18
`define DIST_CODE19    5'd19
`define DIST_CODE20    5'd20
`define DIST_CODE21    5'd21
`define DIST_CODE22    5'd22
`define DIST_CODE23    5'd23
`define DIST_CODE24    5'd24
`define DIST_CODE25    5'd25
`define DIST_CODE26    5'd26
`define DIST_CODE27    5'd27
`define DIST_CODE28    5'd28
`define DIST_CODE29    5'd29

`endif